

module ProgramCounter(
    clk_i,
	rst_i,
	pc_write_i,
	pc_in_i,
	pc_out_o
	);
     
//I/O ports
input           clk_i;
input	        rst_i;
input           pc_write_i;
input  [32-1:0] pc_in_i;
output [32-1:0] pc_out_o;
 
//Internal Signals
logic    [32-1:0] pc_out_o;
 
//Parameter

    
//Main function
always_ff @(posedge clk_i) begin
    if(~rst_i)
	    pc_out_o <= 0;
	else if(pc_write_i)
	    pc_out_o <= pc_in_i;
	else
	    pc_out_o = pc_out_o - 4;
end

endmodule



                    
                    
